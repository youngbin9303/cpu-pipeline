module shift_register
(
	input clk,
	input load,
	input datain,
	output logic dataout
);
